module control(output [8:0] control_bus, input [31:26] op);



endmodule